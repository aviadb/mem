*Model Description
.param temp=27
.param supl = 1.8V

*Including sky130 device models
.lib "sky130_fd_pr/models/sky130.lib.spice" tt


Vdd vdd 0 {supl}

* transistors
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 w=1.05 l=.15 m=1
XM2 out in 0 0 sky130_fd_pr__nfet_01v8 w=.42 l=.15 m=1


Cload out 0 1fF

* input
Vin in 0 1.8

.op
.dc Vin 0 1.8 0.02

.control
run 
display
setplot
setplot dc1
display
plot out vs in
.endc

.end